module instr_mem(
    input logic     A.
    output logic    RD
);