module sign_extend(
    input logic     ImmSrc,
    input logic     instr,
    output logic    ImmOp
)