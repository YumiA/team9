module ALU #(

) (

)

endmodule